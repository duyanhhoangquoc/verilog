module encode3to8(sel1, sel2, sel3, out);
input sel1, sel2, sel3;
output reg [7:0] out;

always @(sel1, sel2, sel3) begin
    case ({sel1, sel2, sel3})
        3'b000: out = 8'b10000000; //if ((sel1, sel2, sel3) == 3'b00)
        3'b001: out = 8'b01000000;
        3'b010: out = 8'b00100000;
        3'b011: out = 8'b00010000;
        3'b100: out = 8'b00001000;
        3'b101: out = 8'b00000100;
        3'b110: out = 8'b00000010;
        3'b111: out = 8'b00000001;
        default: out = 8'b00000000;
    endcase
end
endmodule